`timescale 1ns/1ns
module cmos_capture_raw_gray
#(
	parameter	CMOS_FRAME_WAITCNT	=	4'd10  //等待数据稳定所需要的帧数
															
)
(
	//global clock
	input		clk_cmos,			           //锁相环分频时钟
	input		rst_n,				           //复位信号，低有效

	//CMOS Sensor Interface
	input		cmos_pclk,			           //摄像头输入时钟
	output		cmos_xclk,			           //摄像头驱动时钟
	input		cmos_vsync,			           //摄像头场信号
	input		cmos_href,					   //摄像头行信号
	input [7:0]	cmos_data,					   //摄像头数据
	
	//CMOS SYNC Data output
    output		cmos_frame_vsync,			   //摄像头场有效信号
    output		cmos_frame_href,			   //摄像头行有效信号
    output[7:0]wr_data,			           //摄像头有效数据	
    output		cmos_frame_clken,			   //摄像头数据有效使能
	
	//user interface
	output reg[7:0]	cmos_fps_rate				   //摄像头帧率
);

//parameter define   
localparam	DELAY_TOP = 2 * 24_000000;	//2s delay

//reg define
reg	[27:0]	delay_cnt;
reg		    frame_sync_flag;  //判断有效帧 （10帧后）
reg	[3:0]	cmos_fps_cnt;
reg	[1:0]	cmos_vsync_r, cmos_href_r; //低位是当前 clock 高位是延时一位的clk
reg	[7:0]	cmos_data_r0, cmos_data_r1;
reg	[8:0]	cmos_fps_cnt2;

//wire define
wire        cmos_vsync_end;
wire        delay_2s;
wire [7:0]  cmos_frame_data;

//*****************************************************
//**                    main code
//*****************************************************   

assign	cmos_vsync_end 		= 	(cmos_vsync_r[1] & ~cmos_vsync_r[0]) ? 1'b1 : 1'b0;	
assign	cmos_xclk = clk_cmos;	//24MHz CMOS XCLK output
assign	cmos_frame_clken = frame_sync_flag  ? cmos_href_r[1] : 1'b0;
assign	cmos_frame_vsync = frame_sync_flag  ? cmos_vsync_r[1] : 1'b0;//DFF 2 clocks 输出的同步信号是输入的延时
assign	cmos_frame_href  = frame_sync_flag ? cmos_href_r[1] : 1'b0;	//DFF 2 clocks  
assign	cmos_frame_data	 = frame_sync_flag  ? cmos_data_r1 : 8'd0;	//DFF 2 clocks
assign	delay_2s = (delay_cnt == DELAY_TOP - 1'b1) ? 1'b1 : 1'b0;
assign	wr_data = cmos_frame_data;
//assign  wr_data = {cmos_frame_data[7:3],cmos_frame_data[7:2],cmos_frame_data[7:3]};

//信号延时
always@(posedge cmos_pclk or negedge rst_n)begin
	if(!rst_n)
		begin
		cmos_vsync_r <= 0;
		cmos_href_r <= 0;
		cmos_data_r0 <= 8'd0;
		cmos_data_r1 <= 8'd0;
		end
	else
		begin
		cmos_vsync_r <= {cmos_vsync_r[0], cmos_vsync};
		cmos_href_r <= {cmos_href_r[0], cmos_href};
		cmos_data_r0 <= cmos_data;
		cmos_data_r1 <= cmos_data_r0;
//		{cmos_data_r1, cmos_data_r0} <= {cmos_data_r0, cmos_data};
		end
end

//Wait for Sensor output Data valid 10 Frame of OmniVision
always@(posedge cmos_pclk or negedge rst_n)begin
	if(!rst_n)
		cmos_fps_cnt <= 0;
	else	//Wait until cmos init complete
		begin
		if(cmos_fps_cnt < CMOS_FRAME_WAITCNT)	
			cmos_fps_cnt <= cmos_vsync_end ? cmos_fps_cnt + 1'b1 : cmos_fps_cnt;
		else
			cmos_fps_cnt <= CMOS_FRAME_WAITCNT;  //帧页面记数
		end
end

//Come ture frame synchronization to ignore error frame or has not capture when vsync begin
always@(posedge cmos_pclk or negedge rst_n)begin
	if(!rst_n)
		frame_sync_flag <= 0;
	else if(cmos_fps_cnt == CMOS_FRAME_WAITCNT && cmos_vsync_end == 1)
		frame_sync_flag <= 1;
	else
		frame_sync_flag <= frame_sync_flag;
end

//Delay 2s for cmos fps counter
always@(posedge cmos_pclk or negedge rst_n)begin
	if(!rst_n)
		delay_cnt <= 0;
	else if(delay_cnt < DELAY_TOP - 1'b1)
		delay_cnt <= delay_cnt + 1'b1;
	else
		delay_cnt <= 0;
end

//cmos image output rate counter
always@(posedge cmos_pclk or negedge rst_n)begin
	if(!rst_n)
		begin
		cmos_fps_cnt2 <= 0;
		cmos_fps_rate <= 0;
		end
	else if(delay_2s == 1'b0)	//time is not reached
		begin
		cmos_fps_cnt2 <= cmos_vsync_end ? cmos_fps_cnt2 + 1'b1 : cmos_fps_cnt2;
		cmos_fps_rate <= cmos_fps_rate;
		end
	else	//time up
		begin
		cmos_fps_cnt2 <= 0;
		cmos_fps_rate <= cmos_fps_cnt2[8:1];	//divide by 2
		end
end

endmodule
